module ADC(

); 

endmodule 